BZh91AY&SY��	� i߀Py����߰����P~t�ٝ�  i(Ѧ�Pi����@h��J�I�Q��6�z� d4�ѐ@Jh��1 �di�G�ɠ��� c��4�	��0#F�` @�$�2	�!4�H�O��xP4�3D�?r%����?ʍ�%�?�������_�:���IT%Ra��mBxTb�^�*5a�7n�	0�
�Q��JC;&�]���)m��MV�[�lb���y�]�L�+$�[�k'[�-����m��_M����d+"�:����C�6Y<�Y�RKT]e�T���Nk`�٩u�l^�)J���:�k�4�8��Qe`l�rIC	��$�C��Z.4��"{����@�Yv�ɤ���ɛ62��
O��I�OCb�Z��Q�Mτ�M*k����j��ի�ਭ�1�9<�6�m���)�
��"-Nw���d��Yi-���f��b$�)�����Cm�4@H���c�n-�#�㠒%�Q��[�}H��k.H�<�U=��'*|��Zܻ�%8=K�����Y��azI���פ5�j�=�{꺤��,�^��6�+uSn�U'���k�ò��Ӓ�l4c�ɲڕf;�4k���9}&+H�B��p����xCjg��j�f�3�V{e��+�W���(����iA��>/���c(�u˳�Cv�r�vn8���'բ�i)i�wu?6�
2�]�)��0��)�Q���-n\*��sj:ԩ7㩱�5�����D�^<������Y;�%6�M�O��p�OvF�4lczT���V9"�¶-�f�i��o�睡|6-��8Q]W�e"�f#�s�.���/t��p���'���>i�oquI�X,���7�:����)�ܓ�x�J�7�i��4T�ʪE�q��t�y����;Z7z�;7HŰSt��T��έ*�v���;:7~ڰ�}�Ne�p��gǥ�����L;v8b����3��N&CQ0%�n�~��e�ĝ�u7�7����-�4�tK�F��߂�R���&�a����"�(HMW� 